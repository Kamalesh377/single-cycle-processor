:(
  
